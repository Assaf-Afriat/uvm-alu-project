
// UVM Environment
// Top-level verification component.

class alu_env extends uvm_env;
    `uvm_component_utils(alu_env)

    alu_agent      agent;
    alu_scoreboard scoreboard;

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        agent      = alu_agent::type_id::create("agent", this);
        scoreboard = alu_scoreboard::type_id::create("scoreboard", this);
    endfunction

    function void connect_phase(uvm_phase phase);
        // Connect Monitor -> Scoreboard (2 channels)
        agent.monitor.req_port.connect(scoreboard.req_export);
        agent.monitor.resp_port.connect(scoreboard.resp_export);
    endfunction

endclass
